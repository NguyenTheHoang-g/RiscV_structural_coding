module control_logic(
input logic [10:0] address,
output logic [11:0] ctrl_signal);

	 logic [11:0] rom[0:2047];
	 initial begin
	 rom[11'b01100_000_0_0_0] = 12'b0_1_0_0_0_0000_01_0;  // ADD
	 rom[11'b01100_000_0_0_1] = 12'b0_1_0_0_0_0000_01_0;  
	 rom[11'b01100_000_0_1_0] = 12'b0_1_0_0_0_0000_01_0;  
	 rom[11'b01100_000_0_1_1] = 12'b0_1_0_0_0_0000_01_0;  
	 //
	 rom[11'b01100_001_0_0_0] = 12'b0_1_0_0_0_0001_01_0;  // SLL
	 rom[11'b01100_001_0_0_1] = 12'b0_1_0_0_0_0001_01_0;  
	 rom[11'b01100_001_0_1_0] = 12'b0_1_0_0_0_0001_01_0;  
	 rom[11'b01100_001_0_1_1] = 12'b0_1_0_0_0_0001_01_0;  
	 //
	 rom[11'b01100_011_0_0_0] = 12'b0_1_0_0_0_0011_01_0;  // SLU
	 rom[11'b01100_011_0_0_1] = 12'b0_1_0_0_0_0011_01_0;  
	 rom[11'b01100_011_0_1_0] = 12'b0_1_0_0_0_0011_01_0;  
	 rom[11'b01100_011_0_1_1] = 12'b0_1_0_0_0_0011_01_0;
	 //
	 rom[11'b01100_100_0_0_0] = 12'b0_1_0_0_0_0100_01_0;  // XOR
	 rom[11'b01100_100_0_0_1] = 12'b0_1_0_0_0_0100_01_0;  
	 rom[11'b01100_100_0_1_0] = 12'b0_1_0_0_0_0100_01_0;  
	 rom[11'b01100_100_0_1_1] = 12'b0_1_0_0_0_0100_01_0;
	 //
	 rom[11'b01100_010_0_0_0] = 12'b0_1_0_0_0_0010_01_0;  // SLT
	 rom[11'b01100_010_0_0_1] = 12'b0_1_0_0_0_0010_01_0;  
	 rom[11'b01100_010_0_1_0] = 12'b0_1_0_0_0_0010_01_0;  
	 rom[11'b01100_010_0_1_1] = 12'b0_1_0_0_0_0010_01_0;  
	 //
	 rom[11'b01100_101_0_0_0] = 12'b0_1_0_0_0_0101_01_0;  // SLR
	 rom[11'b01100_101_0_0_1] = 12'b0_1_0_0_0_0101_01_0;  
	 rom[11'b01100_101_0_1_0] = 12'b0_1_0_0_0_0101_01_0;  
	 rom[11'b01100_101_0_1_1] = 12'b0_1_0_0_0_0101_01_0;
	 //
	 rom[11'b01100_110_0_0_0] = 12'b0_1_0_0_0_0110_01_0;  // OR
	 rom[11'b01100_110_0_0_1] = 12'b0_1_0_0_0_0110_01_0;  
	 rom[11'b01100_110_0_1_0] = 12'b0_1_0_0_0_0110_01_0;  
	 rom[11'b01100_110_0_1_1] = 12'b0_1_0_0_0_0110_01_0;
	 //
	 rom[11'b01100_111_0_0_0] = 12'b0_1_0_0_0_0111_01_0;  // AND
	 rom[11'b01100_111_0_0_1] = 12'b0_1_0_0_0_0111_01_0;  
	 rom[11'b01100_111_0_1_0] = 12'b0_1_0_0_0_0111_01_0;  
	 rom[11'b01100_111_0_1_1] = 12'b0_1_0_0_0_0111_01_0;
    //
	 rom[11'b01100_000_1_0_0] = 12'b0_1_0_0_0_1000_01_0;  // ADD
	 rom[11'b01100_000_1_0_1] = 12'b0_1_0_0_0_1000_01_0;  
	 rom[11'b01100_000_1_1_0] = 12'b0_1_0_0_0_1000_01_0;  
	 rom[11'b01100_000_1_1_1] = 12'b0_1_0_0_0_1000_01_0; 
	 //
	 rom[11'b01100_101_1_0_0] = 12'b0_1_0_0_0_1101_01_0;  // SLR
	 rom[11'b01100_101_1_0_1] = 12'b0_1_0_0_0_1101_01_0;  
	 rom[11'b01100_101_1_1_0] = 12'b0_1_0_0_0_1101_01_0;  
	 rom[11'b01100_101_1_1_1] = 12'b0_1_0_0_0_1101_01_0;
	 //
	    // ADDI
    rom[11'b00100_000_0_0_0] = 12'b0_1_0_0_1_0000_01_0;
    rom[11'b00100_000_0_0_1] = 12'b0_1_0_0_1_0000_01_0;
    rom[11'b00100_000_0_1_0] = 12'b0_1_0_0_1_0000_01_0;
    rom[11'b00100_000_0_1_1] = 12'b0_1_0_0_1_0000_01_0;
    //

    // XORI
    rom[11'b00100_100_0_0_0] = 12'b0_1_0_0_1_0100_01_0;
    rom[11'b00100_100_0_0_1] = 12'b0_1_0_0_1_0100_01_0;
    rom[11'b00100_100_0_1_0] = 12'b0_1_0_0_1_0100_01_0;
    rom[11'b00100_100_0_1_1] = 12'b0_1_0_0_1_0100_01_0;
    //

    // ORI
    rom[11'b00100_110_0_0_0] = 12'b0_1_0_0_1_0110_01_0;
    rom[11'b00100_110_0_0_1] = 12'b0_1_0_0_1_0110_01_0;
    rom[11'b00100_110_0_1_0] = 12'b0_1_0_0_1_0110_01_0;
    rom[11'b00100_110_0_1_1] = 12'b0_1_0_0_1_0110_01_0;
    //

    // ANDI
    rom[11'b00100_111_0_0_0] = 12'b0_1_0_0_1_0111_01_0;
    rom[11'b00100_111_0_0_1] = 12'b0_1_0_0_1_0111_01_0;
    rom[11'b00100_111_0_1_0] = 12'b0_1_0_0_1_0111_01_0;
    rom[11'b00100_111_0_1_1] = 12'b0_1_0_0_1_0111_01_0;
    //

    // SLLI
    rom[11'b00100_001_0_0_0] = 12'b0_1_0_0_1_0001_01_0;
    rom[11'b00100_001_0_0_1] = 12'b0_1_0_0_1_0001_01_0;
    rom[11'b00100_001_0_1_0] = 12'b0_1_0_0_1_0001_01_0;
    rom[11'b00100_001_0_1_1] = 12'b0_1_0_0_1_0001_01_0;
    //

    // SRLI
    rom[11'b00100_101_0_0_0] = 12'b0_1_0_0_1_0101_01_0;
    rom[11'b00100_101_0_0_1] = 12'b0_1_0_0_1_0101_01_0;
    rom[11'b00100_101_0_1_0] = 12'b0_1_0_0_1_0101_01_0;
    rom[11'b00100_101_0_1_1] = 12'b0_1_0_0_1_0101_01_0;
    //

    // SRAI
    rom[11'b00100_101_1_0_0] = 12'b0_1_0_0_1_1101_01_0;
    rom[11'b00100_101_1_0_1] = 12'b0_1_0_0_1_1101_01_0;
    rom[11'b00100_101_1_1_0] = 12'b0_1_0_0_1_1101_01_0;
    rom[11'b00100_101_1_1_1] = 12'b0_1_0_0_1_1101_01_0;
    //

    // SLTI
    rom[11'b00100_010_0_0_0] = 12'b0_1_0_0_1_0100_01_0;
    rom[11'b00100_010_0_0_1] = 12'b0_1_0_0_1_0100_01_0;
    rom[11'b00100_010_0_1_0] = 12'b0_1_0_0_1_0100_01_0;
    rom[11'b00100_010_0_1_1] = 12'b0_1_0_0_1_0100_01_0;
    //

    // SLTIU
    rom[11'b00100_011_0_0_0] = 12'b0_1_0_0_1_0011_01_0;
    rom[11'b00100_011_0_0_1] = 12'b0_1_0_0_1_0011_01_0;
    rom[11'b00100_011_0_1_0] = 12'b0_1_0_0_1_0011_01_0;
    rom[11'b00100_011_0_1_1] = 12'b0_1_0_0_1_0011_01_0;
    //
	 // LH
	 rom[11'b00000_000_0_0_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_000_0_0_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_000_0_1_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_000_0_1_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_000_1_0_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_000_1_0_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_000_1_1_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_000_1_1_1] = 12'b1_1_0_0_1_0000_10_0;
    // 
	 // LW
	 rom[11'b00000_001_0_0_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_001_0_0_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_001_0_1_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_001_0_1_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_001_1_0_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_001_1_0_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_001_1_1_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_001_1_1_1] = 12'b1_1_0_0_1_0000_10_0;
	 //
	 // LBU
	 rom[11'b00000_100_0_0_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_100_0_0_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_100_0_1_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_100_0_1_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_100_1_0_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_100_1_0_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_100_1_1_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_100_1_1_1] = 12'b1_1_0_0_1_0000_10_0;
	 //
	 //LHU
	 rom[11'b00000_101_0_0_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_101_0_0_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_101_0_1_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_101_0_1_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_101_1_0_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_101_1_0_1] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_101_1_1_0] = 12'b1_1_0_0_1_0000_10_0;
	 rom[11'b00000_101_1_1_1] = 12'b1_1_0_0_1_0000_10_0;
	 //
	 //SB
	 rom[11'b01000_000_0_0_0] = 12'b0_0_0_0_1_0000_00_1;
	 rom[11'b01000_000_0_0_1] = 12'b0_0_0_0_1_0000_01_1;
	 rom[11'b01000_000_0_1_0] = 12'b0_0_0_0_1_0000_10_1;
	 rom[11'b01000_000_0_1_1] = 12'b0_0_0_0_1_0000_11_1;
	 rom[11'b01000_000_1_0_0] = 12'b0_0_1_0_1_0000_00_1;
	 rom[11'b01000_000_1_0_1] = 12'b0_0_1_0_1_0000_01_1;
	 rom[11'b01000_000_1_1_0] = 12'b0_0_1_0_1_0000_10_1;
	 rom[11'b01000_000_1_1_1] = 12'b0_0_1_0_1_0000_11_1;
	 //
	 //SH
	 rom[11'b01000_001_0_0_0] = 12'b0_0_0_0_1_0000_00_1;
	 rom[11'b01000_001_0_0_1] = 12'b0_0_0_0_1_0000_01_1;
	 rom[11'b01000_001_0_1_0] = 12'b0_0_0_0_1_0000_10_1;
	 rom[11'b01000_001_0_1_1] = 12'b0_0_0_0_1_0000_11_1;
	 rom[11'b01000_001_1_0_0] = 12'b0_0_1_0_1_0000_00_1;
	 rom[11'b01000_001_1_0_1] = 12'b0_0_1_0_1_0000_01_1;
	 rom[11'b01000_001_1_1_0] = 12'b0_0_1_0_1_0000_10_1;
	 rom[11'b01000_001_1_1_1] = 12'b0_0_1_0_1_0000_11_1;
	 //
	 //SW
	 rom[11'b01000_010_0_0_0] = 12'b0_0_0_0_1_0000_00_1;
	 rom[11'b01000_010_0_0_1] = 12'b0_0_0_0_1_0000_01_1;
	 rom[11'b01000_010_0_1_0] = 12'b0_0_0_0_1_0000_10_1;
	 rom[11'b01000_010_0_1_1] = 12'b0_0_0_0_1_0000_11_1;
	 rom[11'b01000_010_1_0_0] = 12'b0_0_1_0_1_0000_00_1;
	 rom[11'b01000_010_1_0_1] = 12'b0_0_1_0_1_0000_01_1;
	 rom[11'b01000_010_1_1_0] = 12'b0_0_1_0_1_0000_10_1;
	 rom[11'b01000_010_1_1_1] = 12'b0_0_1_0_1_0000_11_1;
	 //
	 //BEQ
	 rom[11'b11000_000_0_0_1] = 12'b1_0_0_1_1_0000_01_0;
	 rom[11'b11000_000_1_0_1] = 12'b1_0_0_1_1_0000_01_0;
	
  	 rom[11'b11000_000_0_0_0] = 12'b0_0_0_1_1_0000_01_0;
	 rom[11'b11000_000_0_1_0] = 12'b0_0_0_1_1_0000_01_0;
	 rom[11'b11000_000_1_0_0] = 12'b0_0_0_1_1_0000_01_0;
	 rom[11'b11000_000_1_1_0] = 12'b0_0_0_1_1_0000_01_0;
	 //
	 //BNE
	 rom[11'b11000_001_0_0_0] = 12'b1_0_0_1_1_0000_01_0;
	 rom[11'b11000_001_0_1_0] = 12'b1_0_0_1_1_0000_01_0;
	 rom[11'b11000_001_1_0_0] = 12'b1_0_0_1_1_0000_01_0;
	 rom[11'b11000_001_1_1_0] = 12'b1_0_0_1_1_0000_01_0;
	 
	 rom[11'b11000_001_0_0_1] = 12'b0_0_0_1_1_0000_01_0;
	 rom[11'b11000_001_0_1_1] = 12'b0_0_0_1_1_0000_01_0;
	 rom[11'b11000_001_1_0_1] = 12'b0_0_0_1_1_0000_01_0;
	 rom[11'b11000_001_1_1_1] = 12'b0_0_0_1_1_0000_01_0;
	 //
	 //BLT
	 rom[11'b11000_100_0_1_0] = 12'b1_0_0_1_1_0000_01_0;
	 rom[11'b11000_100_1_1_0] = 12'b1_0_0_1_1_0000_01_0;
	 
	 rom[11'b11000_100_0_0_0] = 12'b0_0_0_1_1_0000_01_0;
	 rom[11'b11000_100_0_0_1] = 12'b0_0_0_1_1_0000_01_0;
	 rom[11'b11000_100_1_0_0] = 12'b0_0_0_1_1_0000_01_0;
	 rom[11'b11000_100_1_0_1] = 12'b0_0_0_1_1_0000_01_0;
	 //
	 //BGE
	 rom[11'b11000_101_0_0_1] = 12'b1_0_0_1_1_0000_01_0;
	 rom[11'b11000_101_1_0_1] = 12'b1_0_0_1_1_0000_01_0;
	 
	 rom[11'b11000_101_0_1_0] = 12'b0_0_0_1_1_0000_01_0;
	 rom[11'b11000_101_1_1_0] = 12'b0_0_0_1_1_0000_01_0;
	 //
	 //BLTU
	 rom[11'b11000_110_0_1_0] = 12'b1_0_1_1_1_0000_01_0;
	 rom[11'b11000_110_1_1_0] = 12'b1_0_1_1_1_0000_01_0;
	 
	 rom[11'b11000_110_0_0_0] = 12'b0_0_1_1_1_0000_01_0;
	 rom[11'b11000_110_0_0_1] = 12'b0_0_1_1_1_0000_01_0;
	 rom[11'b11000_110_1_0_0] = 12'b0_0_1_1_1_0000_01_0;
	 rom[11'b11000_110_1_0_1] = 12'b0_0_1_1_1_0000_01_0;
	 //
	 //BGEU
	 rom[11'b11000_111_0_0_1] = 12'b1_0_1_1_1_0000_01_0;
	 rom[11'b11000_111_1_0_1] = 12'b1_0_1_1_1_0000_01_0;
	 
	 rom[11'b11000_111_0_0_1] = 12'b0_0_1_1_1_0000_01_0;
	 rom[11'b11000_111_1_0_1] = 12'b0_0_1_1_1_0000_01_0;
	 //
	 //JAL
	 rom[11'b11011_000_0_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_000_0_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_000_0_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_000_0_1_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_000_1_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_000_1_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_000_1_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_000_1_1_1] = 12'b1_1_0_1_1_0000_00_0;

	rom[11'b11011_001_0_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_001_0_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_001_0_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_001_0_1_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_001_1_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_001_1_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_001_1_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_001_1_1_1] = 12'b1_1_0_1_1_0000_00_0;

	rom[11'b11011_010_0_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_010_0_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_010_0_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_010_0_1_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_010_1_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_010_1_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_010_1_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_010_1_1_1] = 12'b1_1_0_1_1_0000_00_0;

	rom[11'b11011_011_0_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_011_0_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_011_0_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_011_0_1_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_011_1_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_011_1_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_011_1_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_011_1_1_1] = 12'b1_1_0_1_1_0000_00_0;

	rom[11'b11011_100_0_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_100_0_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_100_0_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_100_0_1_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_100_1_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_100_1_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_100_1_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_100_1_1_1] = 12'b1_1_0_1_1_0000_00_0;

	rom[11'b11011_101_0_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_101_0_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_101_0_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_101_0_1_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_101_1_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_101_1_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_101_1_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_101_1_1_1] = 12'b1_1_0_1_1_0000_00_0;

	rom[11'b11011_110_0_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_110_0_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_110_0_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_110_0_1_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_110_1_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_110_1_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_110_1_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_110_1_1_1] = 12'b1_1_0_1_1_0000_00_0;

	rom[11'b11011_111_0_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_111_0_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_111_0_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_111_0_1_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_111_1_0_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_111_1_0_1] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_111_1_1_0] = 12'b1_1_0_1_1_0000_00_0;
	rom[11'b11011_111_1_1_1] = 12'b1_1_0_1_1_0000_00_0;
	//
	//JALR
	rom[11'b11001_000_0_0_0] = 12'b1_1_0_0_1_0000_00_0;
	rom[11'b11001_000_0_0_1] = 12'b1_1_0_0_1_0000_00_0;
	rom[11'b11001_000_0_1_0] = 12'b1_1_0_0_1_0000_00_0;
	rom[11'b11001_000_0_1_1] = 12'b1_1_0_0_1_0000_00_0;
	rom[11'b11001_000_1_0_0] = 12'b1_1_0_0_1_0000_00_0;
	rom[11'b11001_000_1_0_1] = 12'b1_1_0_0_1_0000_00_0;
	rom[11'b11001_000_1_1_0] = 12'b1_1_0_0_1_0000_00_0;
	rom[11'b11001_000_1_1_1] = 12'b1_1_0_0_1_0000_00_0;
	//
	//LUI
	rom[11'b01101_000_0_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_000_0_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_000_0_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_000_0_1_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_000_1_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_000_1_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_000_1_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_000_1_1_1] = 12'b0_1_0_0_1_0001_01_0;

	rom[11'b01101_001_0_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_001_0_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_001_0_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_001_0_1_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_001_1_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_001_1_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_001_1_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_001_1_1_1] = 12'b0_1_0_0_1_0001_01_0;

	rom[11'b01101_010_0_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_010_0_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_010_0_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_010_0_1_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_010_1_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_010_1_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_010_1_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_010_1_1_1] = 12'b0_1_0_0_1_0001_01_0;

	rom[11'b01101_011_0_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_011_0_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_011_0_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_011_0_1_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_011_1_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_011_1_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_011_1_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_011_1_1_1] = 12'b0_1_0_0_1_0001_01_0;

	rom[11'b01101_100_0_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_100_0_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_100_0_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_100_0_1_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_100_1_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_100_1_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_100_1_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_100_1_1_1] = 12'b0_1_0_0_1_0001_01_0;

	rom[11'b01101_101_0_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_101_0_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_101_0_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_101_0_1_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_101_1_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_101_1_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_101_1_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_101_1_1_1] = 12'b0_1_0_0_1_0001_01_0;

	rom[11'b01101_110_0_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_110_0_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_110_0_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_110_0_1_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_110_1_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_110_1_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_110_1_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_110_1_1_1] = 12'b0_1_0_0_1_0001_01_0;

	rom[11'b01101_111_0_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_111_0_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_111_0_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_111_0_1_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_111_1_0_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_111_1_0_1] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_111_1_1_0] = 12'b0_1_0_0_1_0001_01_0;
	rom[11'b01101_111_1_1_1] = 12'b0_1_0_0_1_0001_01_0;
	//
	//AUIPC
	rom[11'b00101_000_0_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_000_0_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_000_0_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_000_0_1_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_000_1_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_000_1_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_000_1_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_000_1_1_1] = 12'b0_1_0_1_1_0000_01_0;

	rom[11'b00101_001_0_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_001_0_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_001_0_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_001_0_1_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_001_1_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_001_1_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_001_1_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_001_1_1_1] = 12'b0_1_0_1_1_0000_01_0;

	rom[11'b00101_010_0_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_010_0_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_010_0_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_010_0_1_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_010_1_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_010_1_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_010_1_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_010_1_1_1] = 12'b0_1_0_1_1_0000_01_0;

	rom[11'b00101_011_0_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_011_0_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_011_0_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_011_0_1_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_011_1_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_011_1_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_011_1_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_011_1_1_1] = 12'b0_1_0_1_1_0000_01_0;

	rom[11'b00101_100_0_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_100_0_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_100_0_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_100_0_1_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_100_1_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_100_1_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_100_1_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_100_1_1_1] = 12'b0_1_0_1_1_0000_01_0;

	rom[11'b00101_101_0_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_101_0_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_101_0_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_101_0_1_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_101_1_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_101_1_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_101_1_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_101_1_1_1] = 12'b0_1_0_1_1_0000_01_0;

	rom[11'b00101_110_0_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_110_0_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_110_0_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_110_0_1_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_110_1_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_110_1_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_110_1_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_110_1_1_1] = 12'b0_1_0_1_1_0000_01_0;

	rom[11'b00101_111_0_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_111_0_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_111_0_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_111_0_1_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_111_1_0_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_111_1_0_1] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_111_1_1_0] = 12'b0_1_0_1_1_0000_01_0;
	rom[11'b00101_111_1_1_1] = 12'b0_1_0_1_1_0000_01_0;
	
	end
	
assign ctrl_signal= rom[address];
endmodule

	

	

	 
	 
	 
	 
	 
	 

	 


	 
