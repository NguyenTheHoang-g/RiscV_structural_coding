module Instruction_mem(
input logic clk, rst,
input logic [31:0] read_addr,
output logic [31:0] instruction_out);

endmodule